module axi_spi_slave #(

)(

);

endmodule
